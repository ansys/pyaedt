*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
C1 2 0 1.967E-12
Ln1L2 2000 2 1E-09
L2 2000 3001 1.288E-08
Ln2L2 3001 3 1E-09
C3 3 0 6.366E-12
Ln1L4 3000 3 1E-09
L4 3000 4001 1.288E-08
Ln2L4 4001 4 1E-09
C5 4 0 1.967E-12
R6 4 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(4) -80 0
.PLOT AC VP(4) -200 200
.PLOT AC VG(4) 0 9E-10
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(4) -0.1 0.6
.END
