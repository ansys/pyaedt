*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
L1 2 3 4.918E-09
C2 3 0 5.15E-12
L3 3 4 1.592E-08
C4 4 0 5.15E-12
L5 4 5 4.918E-09
R6 5 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(5) -80 0
.PLOT AC VP(5) -200 200
.PLOT AC VG(5) 0 9E-10
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(5) 0 0.6
.END
