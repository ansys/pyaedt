*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
*
* Dummy Resistors Required For Spice
* Have Been Added to Net List.
*
C1 2 0 2.29E-13
C2 2 3 4.93E-12
C3 3 0 1.162E-12
L5 3 4 3.706E-09
C6 4 5 2.586E-11
Rq6 4 5 5E+10
C4 3 5 5.248E-12
L7 5 6 8.386E-10
C7 6 0 1.652E-11
C8 5 6 3.079E-11
C10 5 7 2.923E-13
Rq10 5 7 5E+10
L11 7 8 7.329E-08
C9 5 8 3.421E-12
L12 8 9 1.405E-07
C12 9 0 -2.474E-13
C13 8 9 4.788E-13
C14 8 10 -1.186E-11
Rq14 8 10 5E+10
R15 10 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(10) -70 0
.PLOT AC VP(10) -200 200
.PLOT AC VG(10) 0 2E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(10) -0.04 0.08
.END
