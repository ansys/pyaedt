*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
C1 2 0 9.836E-12
L2 2 3 2.476E-09
C3 3 0 2.627E-10
L4 3 4 9.78E-11
C5 4 0 2.04E-08
L6 4 0 1.242E-12
C7 4 5 2.59E-10
L8 5 0 9.641E-11
C9 5 6 1.023E-11
L10 6 0 2.575E-09
R11 6 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(6) -160 0
.PLOT AC VP(6) -200 200
.PLOT AC VG(6) 0 9E-09
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(6) -0.04 0.04
.END
