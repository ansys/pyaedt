*
*Length Units: Meters
*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
Rg 1 2 50
MT1 2 0 Wid=0.001665 Len=0.01084 Er=9.8 Thick=2.54E-06 Height=0.00127
MT2 2 3 Wid=0.001665 Len=0.01697 Er=9.8 Thick=2.54E-06 Height=0.00127
MT3 3 4 Wid=0.001665 Len=0.001888 Er=9.8 Thick=2.54E-06 Height=0.00127
MT4 0 5 3 0 Gap=0.001031 Len=0.02781 Er=9.8 Thick=2.54E-06 Height=0.00127
MT5 5 0 Wid=0.001671 Len=0.02781 Er=9.8 Thick=2.54E-06 Height=0.00127
MT6 5 0 0 6 Gap=0.001726 Len=0.02781 Er=9.8 Thick=2.54E-06 Height=0.00127
MT7 0 6 Wid=0.001749 Len=0.02781 Er=9.8 Thick=2.54E-06 Height=0.00127
MT8 0 7 6 0 Gap=0.001726 Len=0.02781 Er=9.8 Thick=2.54E-06 Height=0.00127
MT9 7 0 Wid=0.001671 Len=0.02781 Er=9.8 Thick=2.54E-06 Height=0.00127
MT10 7 0 0 8 Gap=0.001031 Len=0.02781 Er=9.8 Thick=2.54E-06 Height=0.00127
MT11 0 9 Wid=0.001665 Len=0.01084 Er=9.8 Thick=2.54E-06 Height=0.00127
MT12 9 8 Wid=0.001665 Len=0.01697 Er=9.8 Thick=2.54E-06 Height=0.00127
MT13 8 10 Wid=0.001665 Len=0.001888 Er=9.8 Thick=2.54E-06 Height=0.00127
Rl 9 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(Rl) -80 0
.PLOT AC VP(Rl) -200 200
.PLOT AC VG(Rl) -2E-09 1E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(Rl) -0.04 0.04
.END
