*
*Length Units: Meters
*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
Rg 1 2 50
MXTcoup0 2 3 4 0 Wid=0.0009605 Gap=0.00045 Len=0.02909 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MXTcoup1 4 5 6 0 Wid=0.0006633 Gap=0.0001582 Len=0.02944 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MXTcoup2 6 7 8 0 Wid=0.0005798 Gap=0.0001159 Len=0.02952 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MXTcoup3 8 9 10 0 Wid=0.0006633 Gap=0.0001582 Len=0.02944 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MXTcoup4 10 11 12 0 Wid=0.0009605 Gap=0.00045 Len=0.02909 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
Rl 12 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(Rl) -140 0
.PLOT AC VP(Rl) -200 200
.PLOT AC VG(Rl) -2E-07 5E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(Rl) 0 0.7
.END
