*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 30
C1 2 0 1.865E-12
L2 2 3 4.849E-09
C3 3 0 8.275E-12
L4 3 4 8.956E-09
C5 4 0 8.124E-12
R6 4 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(4) -80 0
.PLOT AC VP(4) -200 200
.PLOT AC VG(4) 0 9E-10
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(4) 0 0.8
.END
