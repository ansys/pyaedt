*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
C1 2 0 6.558E-13
L2 2 3 1.183E-08
C2 3 0 7.587E-13
L3 2 4 1.412E-08
C3 4 0 1.265E-13
L4 2 5 4.292E-09
L5 5 6 4.966E-09
C5 5 6 1.808E-12
L6 6 7 8.281E-10
C6 6 7 2.157E-12
C7 7 0 2.122E-12
L8 7 8 3.657E-09
C8 8 0 2.455E-12
L9 7 9 4.363E-09
C9 9 0 4.095E-13
L10 7 10 4.292E-09
L11 10 11 4.966E-09
C11 10 11 1.808E-12
L12 11 12 8.281E-10
C12 11 12 2.157E-12
C13 12 0 6.558E-13
L14 12 13 1.183E-08
C14 13 0 7.587E-13
L15 12 14 1.412E-08
C15 14 0 1.265E-13
R16 12 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(12) -200 0
.PLOT AC VP(12) -200 200
.PLOT AC VG(12) 0 7E-09
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(12) 0 0.7
.END
