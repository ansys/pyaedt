*
*Length Units: Meters
*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
Rg 1 2 50
MT1S1 2 0 Wid=0.0003175 Len=0.003025 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT1S2 2 6 Wid=0.00508 Len=0.01527 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MTSeg0 2 3 Wid=5E-05 Len=0.06218 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT1S3 3 0 Wid=0.0003175 Len=0.000573 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT1S4 3 9 Wid=0.00508 Len=0.0226 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MTSeg1 3 4 Wid=5E-05 Len=0.06218 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT1S5 4 0 Wid=0.0003175 Len=0.003025 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT1S6 4 12 Wid=0.00508 Len=0.01527 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
Rl 4 0 50
*
* The Following Dummy Resistors May Be Required For Spice.
*
Rstb2 6 0 5E+09
Rstb3 7 0 5E+09
Rseg4 3 0 5E+09
Rstb5 9 0 5E+09
Rstb6 10 0 5E+09
Rstb7 12 0 5E+09
Rstb8 13 0 5E+09
*
* End Dummy Resistors
*
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(Rl) -160 0
.PLOT AC VP(Rl) -200 200
.PLOT AC VG(Rl) -9E-08 1E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(Rl) -0.03 0.03
.END
