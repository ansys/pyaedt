*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
*
* Dummy Resistors Required For Spice
* Have Been Added to Net List.
*
C1 2 0 3.83E-13
C2 2 3 4.123E-12
C3 3 0 9.716E-13
L4 3 4 2.561E-09
C4 3 4 6.314E-12
L5 4 5 6.878E-09
C5 5 0 5.769E-12
C6 4 0 1.075E-11
C7 4 6 3.713E-12
Rq7 4 6 5E+10
L8 6 7 4.542E-10
C8 6 7 4.345E-11
L9 7 8 1.229E-07
C9 8 0 2.644E-13
C10 7 0 -5.118E-13
C11 7 9 -1.186E-11
Rq11 7 9 5E+10
R12 9 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(9) -70 0
.PLOT AC VP(9) -200 200
.PLOT AC VG(9) 0 2E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(9) -0.04 0.08
.END
