*
*Length Units: Meters
*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
Rg 1 2 50
MT1 2 3 Wid=0.0004828 Len=0.02763 Er=9.8 Thick=2.54E-06 Height=0.00127
MT2 2 0 3 4 Gap=0.000635 Len=0.02763 Er=9.8 Thick=2.54E-06 Height=0.00127
MT3 0 4 Wid=0.0004828 Len=0.02763 Er=9.8 Thick=2.54E-06 Height=0.00127
MT4 3 4 Wid=0.0004828 Len=0.000635 Er=9.8 Thick=2.54E-06 Height=0.00127
MT5 0 5 4 0 Gap=0.0008077 Len=0.02763 Er=9.8 Thick=2.54E-06 Height=0.00127
MT6 5 0 Wid=0.001735 Len=0.02763 Er=9.8 Thick=2.54E-06 Height=0.00127
MT7 5 0 0 6 Gap=0.001635 Len=0.02763 Er=9.8 Thick=2.54E-06 Height=0.00127
MT8 0 6 Wid=0.001735 Len=0.02763 Er=9.8 Thick=2.54E-06 Height=0.00127
MT9 0 7 6 0 Gap=0.001635 Len=0.02763 Er=9.8 Thick=2.54E-06 Height=0.00127
MT10 7 0 Wid=0.001735 Len=0.02763 Er=9.8 Thick=2.54E-06 Height=0.00127
MT11 7 0 0 8 Gap=0.0008077 Len=0.02763 Er=9.8 Thick=2.54E-06 Height=0.00127
MT12 0 8 Wid=0.0004828 Len=0.02763 Er=9.8 Thick=2.54E-06 Height=0.00127
MT13 0 9 8 10 Gap=0.000635 Len=0.02763 Er=9.8 Thick=2.54E-06 Height=0.00127
MT14 9 10 Wid=0.0004828 Len=0.02763 Er=9.8 Thick=2.54E-06 Height=0.00127
MT15 8 10 Wid=0.0004828 Len=0.000635 Er=9.8 Thick=2.54E-06 Height=0.00127
Rl 9 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(Rl) -70 0
.PLOT AC VP(Rl) -200 200
.PLOT AC VG(Rl) -3E-08 1E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(Rl) -0.04 0.04
.END
