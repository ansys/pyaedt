*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
*
* Dummy Resistors Required For Spice
* Have Been Added to Net List.
*
C1 2 0 1.886E-12
C2 2 3 6.779E-12
L3 3 4 2.646E-08
C3 4 0 1.5E-12
C4 3 5 2.261E-12
Rq4 3 5 5E+10
L5 5 6 1.297E-07
C5 6 0 2.506E-13
L6 5 7 1.91E-09
C6 5 7 1.034E-11
C7 7 0 1.845E-13
C8 7 8 2.717E-12
Rq8 7 8 5E+10
C9 8 0 1.487E-12
L10 8 9 3.91E-09
C10 8 9 4.135E-12
C11 9 0 1.169E-12
R12 9 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(9) -70 0
.PLOT AC VP(9) -200 200
.PLOT AC VG(9) 0 2E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(9) -0.04 0.08
.END
