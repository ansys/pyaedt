*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
Ln1C1 2 2517 1E-09
C1 2517 2519 1.967E-12
Ln2C1 2519 0 1E-09
L2 2 3 1.288E-08
Ln1C3 3 3517 1E-09
C3 3517 3519 6.366E-12
Ln2C3 3519 0 1E-09
L4 3 4 1.288E-08
Ln1C5 4 4517 1E-09
C5 4517 4519 1.967E-12
Ln2C5 4519 0 1E-09
R6 4 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(4) -140 0
.PLOT AC VP(4) -200 200
.PLOT AC VG(4) 0 1.2E-09
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(4) -0.1 0.6
.END
