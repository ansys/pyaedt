*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
L3 2 3 2.968E-08
C4 3 0 1.302E-11
L5 3 4 2.655E-08
C6 4 0 6.873E-12
L7 4 5 5.937E-09
R8 5 0 50
C9 2 6 8.533E-13
L10 6 0 1.945E-09
C11 6 7 9.541E-13
L12 7 0 3.685E-09
C13 7 8 4.267E-12
R14 8 0 50
C15 2 9 4.12E-13
L16 9 10 6.148E-08
L17 10 0 9.393E-10
C18 10 0 2.697E-11
C19 10 11 4.607E-13
L20 11 12 5.499E-08
L21 12 0 1.779E-09
C22 12 0 1.424E-11
C23 12 13 2.06E-12
L24 13 14 1.23E-08
R25 14 0 50
*
* Compensation Elements
*
L1 2 15 1.86E-08
C1 15 0 3.633E-12
L2 2 16 6.972E-09
C2 16 0 1.362E-12
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(5) VDB(8) VDB(14) -160 0
.PLOT AC VP(5) VP(8) VP(14) -200 200
.PLOT AC VG(5) VG(8) VG(14) -2E-09 9E-09
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(5) V(8) V(14) -0.2 0.7
.END
