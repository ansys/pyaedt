*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
*
* Dummy Resistors Required For Spice
* Have Been Added to Net List.
*
L1 2 0 4.285E-09
C2 2 0 5.911E-12
L3 2 3 7.553E-10
C3 2 3 4.289E-11
L4 3 4 5.905E-10
C4 3 4 3.354E-11
L5 4 5 1.237E-09
Rq5 5 0 5E-08
C6 4 0 2.048E-11
L7 4 6 2.913E-09
C7 4 6 1.225E-11
L8 6 7 2.067E-09
C8 6 7 8.696E-12
L9 7 8 2.068E-09
Rq9 8 0 5E-08
C10 7 0 1.225E-11
R11 7 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(7) -60 0
.PLOT AC VP(7) -200 200
.PLOT AC VG(7) 0 2.5E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(7) -0.04 0.04
.END
