*
*Length Units: Meters
*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
Rg 1 2 50
MT1S1 2 0 Wid=0.00635 Len=0.02672 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MTSeg0 2 3 Wid=5E-05 Len=0.06187 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT1S2 3 0 Wid=0.00635 Len=0.02672 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MTSeg1 3 4 Wid=5E-05 Len=0.06187 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT1S3 4 0 Wid=0.00635 Len=0.02672 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
Rl 4 0 50
*
* The Following Dummy Resistors May Be Required For Spice.
*
Rseg2 3 0 5E+09
*
* End Dummy Resistors
*
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(Rl) -160 0
.PLOT AC VP(Rl) -200 200
.PLOT AC VG(Rl) -1.5E-07 5E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(Rl) -0.09 0.07
.END
