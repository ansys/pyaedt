*
I1 1 0 AC 1 PULSE 0 0.04 0 1.592E-13 0
R0 1 0 50
C1 1 0 1.967E-12
L2 1 2 1.288E-08
C3 2 0 6.366E-12
L4 2 3 1.288E-08
C5 3 0 1.967E-12
R6 3 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC IDB(R6) -80 0
.PLOT AC IP(R6) -200 200
.PLOT AC VG(R6) 0 9E-10
.TRAN  5E-11 1E-08 0
.PLOT TRAN I(R6) 0 0.6
.END
