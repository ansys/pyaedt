*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
*
* Dummy Resistors Required For Spice
* Have Been Added to Net List.
*
L1 2 0 2.575E-09
C2 2 3 1.23E-11
C3 3 0 4.918E-11
L4 3 4 2.575E-09
C5 4 0 1.041E-11
C6 4 5 1.302E-12
Rq6 4 5 5E+10
L7 5 0 2.575E-09
C8 5 0 7.522E-12
C9 5 6 1.302E-12
C10 6 0 1.041E-11
L11 6 7 2.575E-09
C12 7 0 4.918E-11
C13 7 8 1.23E-11
Rq13 7 8 5E+10
L14 8 0 2.575E-09
R15 8 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(8) -160 0
.PLOT AC VP(8) -200 200
.PLOT AC VG(8) 0 9E-09
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(8) -0.04 0.04
.END
