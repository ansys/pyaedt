*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
C1 2 3 1.967E-12
LXcs1 3 0 1E-09
L2 2 4 1.288E-08
C3 4 5 6.366E-12
LXcs3 5 0 1E-09
L4 4 6 1.288E-08
C5 6 7 1.967E-12
LXcs5 7 0 1E-09
R6 6 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(6) -160 0
.PLOT AC VP(6) -200 200
.PLOT AC VG(6) 0 1E-09
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(6) 0 0.6
.END
