*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 98.45
*
* Dummy Resistors Required For Spice
* Have Been Added to Net List.
*
L1 2 0 1.413E-08
C2 2 0 1.455E-12
L3 2 3 1.389E-09
C3 2 3 2.333E-11
C4 3 0 6.44E-13
L5 3 4 9.637E-10
C5 3 4 2.055E-11
L6 4 5 1.841E-09
Rq6 5 0 5E-08
C7 4 0 1.313E-11
L8 4 6 3.952E-09
C8 4 6 9.032E-12
C9 6 0 6.44E-13
L10 6 7 2.251E-09
C10 6 7 7.985E-12
L11 7 8 1.912E-09
Rq11 8 0 5E-08
C12 7 0 1.296E-11
R13 7 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(7) -60 0
.PLOT AC VP(7) -200 200
.PLOT AC VG(7) 0 2.5E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(7) -0.03 0.03
.END
