*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
C1 2 0 1.967E-12
Cn1L2 2 0 1E-09
L2 2 3 1.288E-08
Cn2L2 3 0 1E-09
C3 3 0 6.366E-12
Cn1L4 3 0 1E-09
L4 3 4 1.288E-08
Cn2L4 4 0 1E-09
C5 4 0 1.967E-12
R6 4 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(4) -200 -50
.PLOT AC VP(4) -90 0
.PLOT AC VG(4) 0 3E-11
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(4) -0.1 0.6
.END
