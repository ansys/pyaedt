 5              1
 4              2.033e+10
 3              2.067e+20
 2              1.299e+30
 1              5.044e+39
 0   9.793e+48  9.793e+48
