*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
*
* Dummy Resistors Required For Spice
* Have Been Added to Net List.
*
L1 2 3 2.923E-09
L2 3 0 8.341E-09
L3 3 4 1.034E-08
C3 4 0 1.564E-12
L4 3 5 9.446E-09
C4 3 5 4.201E-12
L5 5 6 9.231E-08
Rq5 6 0 5E-08
L6 5 7 2.175E-08
L7 7 8 1.01E-08
Rq7 8 0 5E-08
L8 7 9 1.086E-07
C8 9 0 1.817E-13
L9 7 10 6.611E-10
C9 7 10 4.918E-11
L10 10 11 -1.28E-09
L11 11 12 -2.966E-08
Rq11 12 0 5E-08
R12 11 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(11) -70 0
.PLOT AC VP(11) -200 200
.PLOT AC VG(11) 0 2E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(11) -0.04 0.08
.END
