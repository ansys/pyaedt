*
*Length Units: Meters
*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
Rg 1 2 50
MT1 2 0 Wid=0.00159 Len=0.005702 Er=9.8 Thick=2.54E-06 Height=0.00127
MT2 2 3 Wid=0.00159 Len=0.007848 Er=9.8 Thick=2.54E-06 Height=0.00127
C2 3 0 4.004E-12
MT3 0 0 3 4 Gap=0.001385 Len=0.01355 Er=9.8 Thick=2.54E-06 Height=0.00127
MT4 0 4 Wid=0.00159 Len=0.01355 Er=9.8 Thick=2.54E-06 Height=0.00127
C4 4 0 3.853E-12
MT5 0 0 4 5 Gap=0.002114 Len=0.01355 Er=9.8 Thick=2.54E-06 Height=0.00127
MT6 0 5 Wid=0.00159 Len=0.01355 Er=9.8 Thick=2.54E-06 Height=0.00127
C6 5 0 3.853E-12
MT7 0 0 5 6 Gap=0.002114 Len=0.01355 Er=9.8 Thick=2.54E-06 Height=0.00127
MT8 0 6 Wid=0.00159 Len=0.01355 Er=9.8 Thick=2.54E-06 Height=0.00127
C8 6 0 3.853E-12
MT9 0 0 6 7 Gap=0.001385 Len=0.01355 Er=9.8 Thick=2.54E-06 Height=0.00127
C9 7 0 4.004E-12
MT10 0 8 Wid=0.00159 Len=0.005702 Er=9.8 Thick=2.54E-06 Height=0.00127
MT11 8 7 Wid=0.00159 Len=0.007848 Er=9.8 Thick=2.54E-06 Height=0.00127
Rl 8 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(Rl) -80 0
.PLOT AC VP(Rl) -200 200
.PLOT AC VG(Rl) 0 1.6E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(Rl) -0.05 0.07
.END
