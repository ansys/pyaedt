*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
C3 2 3 4.12E-13
L4 3 4 6.148E-08
L5 4 0 9.393E-10
C6 4 0 2.697E-11
C7 4 5 4.607E-13
L8 5 6 5.499E-08
L9 6 0 1.779E-09
C10 6 0 1.424E-11
C11 6 7 2.06E-12
L12 7 8 1.23E-08
R13 8 0 50
L14 2 9 2.459E-08
C14 2 9 1.03E-12
L15 9 10 2.348E-09
C15 10 0 1.079E-11
L16 9 11 2.199E-08
C16 9 11 1.152E-12
L17 11 12 4.449E-09
C17 12 0 5.694E-12
L18 11 13 4.918E-09
C18 11 13 5.15E-12
R19 13 0 50
*
* Compensation Elements
*
L1 2 14 1.745E-08
C1 14 0 3.873E-12
L2 2 15 6.54E-09
C2 15 0 1.452E-12
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(8) VDB(13) -200 0
.PLOT AC VP(8) VP(13) -200 200
.PLOT AC VG(8) VG(13) -1E-09 9E-09
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(8) V(13) -0.2 0.7
.END
