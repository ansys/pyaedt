*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
C1 2 0 1.967E-12
L2 2 3 1.288E-08
Rs2 3 4 1
C3 4 0 6.366E-12
L4 4 5 1.288E-08
Rs4 5 6 1
C5 6 0 1.967E-12
R6 6 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(6) -80 0
.PLOT AC VP(6) -200 200
.PLOT AC VG(6) 0 9E-10
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(6) 0 0.6
.END
