
Q7 BUS_N N1781183 N1781293 BUS_N BUS_N N1781293 N1781293 N1781293 STS6NF20V
R379 N1850915 N1850867 10k
D174 OINC VDD_3.3V TMMBAT46
J62 INM-DIAG2_Q3 DIAG1_Q3 SD_Q3 BUS_N CON4
C213 VH_Q1 GND_ISO_Q1 1uF/50V
D142 N1763408 DIAG1_Q2 GREEN
R481 N1803431 VBIAS_DC_CURR definire
C246 CS_Q3 BUS_N 47p/50V
R318 N1721592 N1722018 10k
L200 N1721592 BUS_N 1uH
U48 N1814870 BUS_N N1804444 GND_MEAS_DC DCH010505SN7
V1 N1721592 BUS_N 12
V2 N1814870 0 PULSE(0 10 0 0.1u 0.1u 1.2u 5u)
I1 N1763408 0 1e-3
.param a=50V
.PARAM definire=20
.param a1=50V
.PARAM definire2=20
.param a3=50V
.PARAM definire3=20
.param a4=50V
.PARAM definire4=20
.model CON4 V1
.lib C:\Temp\model.lib
.END
