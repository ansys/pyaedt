*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
*
* Dummy Resistors Required For Spice
* Have Been Added to Net List.
*
L1 2 0 3.08E-09
C2 2 0 9.836E-12
L3 2 3 1.263E-08
L4 3 4 3.08E-09
Rq4 4 0 5E-08
C5 3 0 8.641E-12
C6 3 5 1.589E-12
L7 5 0 1.269E-09
C8 5 0 1.728E-11
C9 5 6 1.589E-12
L10 6 0 3.08E-09
C11 6 0 8.641E-12
L12 6 7 1.263E-08
L13 7 8 3.08E-09
Rq13 8 0 5E-08
C14 7 0 9.836E-12
R15 7 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(7) -160 0
.PLOT AC VP(7) -200 200
.PLOT AC VG(7) 0 9E-09
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(7) -0.04 0.04
.END
