*
*Length Units: Meters
*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
Rg 1 2 50
MTSeg0 2 3 Wid=0.002204 Len=0.02834 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MXTcoup1 4 3 6 5 Wid=0.0009521 Gap=0.0004417 Len=0.0293 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MXTcoup2 7 6 9 8 Wid=0.001061 Gap=0.001016 Len=0.029 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MXTcoup3 10 9 12 11 Wid=0.001061 Gap=0.001016 Len=0.029 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MXTcoup4 13 12 15 14 Wid=0.0009521 Gap=0.0004417 Len=0.0293 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MTSeg5 15 16 Wid=0.002204 Len=0.02834 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
Rl 16 0 50
*
* The Following Dummy Resistors May Be Required For Spice.
*
Rseg6 3 0 5E+09
*
* End Dummy Resistors
*
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(Rl) -160 0
.PLOT AC VP(Rl) -200 200
.PLOT AC VG(Rl) -3E-08 2E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(Rl) -0.06 0.1
.END
