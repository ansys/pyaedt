*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
*
* Dummy Resistors Required For Spice
* Have Been Added to Net List.
*
L1 2 0 4.003E-09
C2 2 0 6.443E-12
L3 2 3 7.648E-10
C3 2 3 4.236E-11
L4 3 4 4.003E-09
Rq4 4 0 5E-08
C5 3 0 4.743E-12
L6 3 5 7.217E-10
C6 3 5 2.744E-11
L7 5 6 4.003E-09
Rq7 6 0 5E-08
C8 5 0 6.711E-12
L9 5 7 3.148E-09
C9 5 7 1.134E-11
L10 7 8 5.758E-09
Rq10 8 0 5E-08
C11 7 0 5.081E-12
L12 7 9 1.851E-09
C12 7 9 9.713E-12
L13 9 10 2.342E-09
Rq13 10 0 5E-08
C14 9 0 1.123E-11
R15 9 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(9) -60 0
.PLOT AC VP(9) -200 200
.PLOT AC VG(9) 0 2.5E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(9) -0.04 0.04
.END
