*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 75
L1 2 0 3.863E-09
C2 2 0 6.499E-12
C3 2 3 3.213E-13
C4 3 0 7.22E-14
L5 3 4 6.438E-08
L6 4 0 7.958E-10
C7 4 0 3.183E-11
C8 4 5 3.935E-13
L9 5 6 6.438E-08
L10 6 0 2.575E-09
C11 6 0 9.836E-12
R12 6 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(6) -160 0
.PLOT AC VP(6) -200 200
.PLOT AC VG(6) 0 9E-09
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(6) -0.03 0.03
.END
