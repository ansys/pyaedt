*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
L3 2 3 3.979E-08
C4 3 0 1.745E-11
L5 3 4 3.559E-08
C6 4 0 9.213E-12
L7 4 5 7.958E-09
R8 5 0 50
C9 2 6 6.366E-13
L10 6 0 1.451E-09
C11 6 7 7.118E-13
L12 7 0 2.749E-09
C13 7 8 3.183E-12
R14 8 0 50
C15 2 9 8.798E-13
L16 9 10 2.879E-08
L17 10 0 2.006E-09
C18 10 0 1.263E-11
C19 10 11 9.836E-13
L20 11 12 2.575E-08
L21 12 0 3.799E-09
C22 12 0 6.667E-12
C23 12 13 4.399E-12
L24 13 14 5.758E-09
R25 14 0 50
*
* Compensation Elements
*
L1 2 15 1.835E-08
C1 15 0 5.521E-12
L2 2 16 4.588E-09
C2 16 0 1.38E-12
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(5) VDB(8) VDB(14) -140 0
.PLOT AC VP(5) VP(8) VP(14) -200 200
.PLOT AC VG(5) VG(8) VG(14) -1E-09 5E-09
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(5) V(8) V(14) -0.2 0.7
.END
