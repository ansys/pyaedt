*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
L3 2 3 3.406E-08
C4 3 0 2.366E-12
L5 3 4 1.693E-08
L2 2 4 1.609E-08
L7 4 5 1.969E-08
C8 5 0 2.523E-12
L9 5 6 7.071E-09
L6 4 6 6.955E-09
R10 6 0 50
*
* Dummy Resistors Required For Spice
* Have Been Added to Net List.
*
C11 2 7 3.1E-12
L12 7 8 1.071E-08
C12 8 0 2.947E-12
C13 7 9 3.118E-12
Rq13 7 9 5E+10
L14 9 10 1.004E-08
C14 10 0 6.135E-12
C15 9 11 1.736E-11
Rq15 9 11 5E+10
R16 11 0 50
*
* Compensation Elements
*
L1 2 12 2.28E-07
C1 12 0 1.111E-13
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(6) VDB(11) -200 0
.PLOT AC VP(6) VP(11) -200 200
.PLOT AC VG(6) VG(11) 0 1.8E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(6) V(11) -0.2 0.7
.END
