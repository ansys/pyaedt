*
*Length Units: Meters
*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
Rg 1 2 50
MXTcoup0 3 2 5 4 Wid=5E-05 Gap=5E-05 Len=0.03147 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MTSeg1 5 6 Wid=5E-05 Len=2.5E-05 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT2S2 6 19 Wid=0.0003175 Len=0.03065 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT1S2 19 17 Wid=0.00508 Len=0.0003439 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT2S3 6 23 Wid=0.0003175 Len=0.01956 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT1S3 23 21 Wid=0.00508 Len=0.0002689 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MTSeg2 6 7 Wid=5E-05 Len=2.5E-05 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MXTcoup3 8 7 10 9 Wid=5E-05 Gap=5E-05 Len=0.03145 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MTSeg4 10 11 Wid=5E-05 Len=2.5E-05 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT2S6 11 29 Wid=0.0003175 Len=0.02845 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT1S6 29 27 Wid=0.00508 Len=0.002097 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT2S7 11 33 Wid=0.0003175 Len=0.0149 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT1S7 33 31 Wid=0.00508 Len=0.00134 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MTSeg5 11 12 Wid=5E-05 Len=2.5E-05 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MXTcoup6 13 12 15 14 Wid=5E-05 Gap=5E-05 Len=0.03147 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
Rl 15 0 50
*
* The Following Dummy Resistors May Be Required For Spice.
*
Rseg7 6 0 5E+09
Rstb8 17 0 5E+09
Rstb9 18 0 5E+09
Rstb10 19 0 5E+09
Rstb11 21 0 5E+09
Rstb12 22 0 5E+09
Rstb13 23 0 5E+09
Rseg14 7 0 5E+09
Rseg15 11 0 5E+09
Rstb16 27 0 5E+09
Rstb17 28 0 5E+09
Rstb18 29 0 5E+09
Rstb19 31 0 5E+09
Rstb20 32 0 5E+09
Rstb21 33 0 5E+09
Rseg22 12 0 5E+09
*
* End Dummy Resistors
*
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(Rl) -120 0
.PLOT AC VP(Rl) -200 200
.PLOT AC VG(Rl) -3E-08 2E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(Rl) -0.04 0.04
.END
