*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
L2 2 3 1.359E-08
C3 3 0 5.96E-12
L4 3 4 1.215E-08
C5 4 0 3.146E-12
L6 4 5 2.717E-09
R7 5 0 50
C8 2 6 1.864E-12
L9 6 0 4.25E-09
C10 6 7 2.084E-12
L11 7 0 8.052E-09
C12 7 8 9.322E-12
R13 8 0 50
*
* Compensation Elements
*
L1 2 9 2.041E-07
C1 9 0 1.241E-13
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(5) VDB(8) -200 0
.PLOT AC VP(5) VP(8) -200 200
.PLOT AC VG(5) VG(8) 0 1.4E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(5) V(8) -0.2 0.7
.END
