*
*Length Units: Meters
*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
Rg 1 2 50
MT1 2 3 Wid=0.00127 Len=0.01137 Er=9.8 Thick=2.54E-06 Height=0.00127
MT2 2 4 Wid=0.00127 Len=0.01424 Er=9.8 Thick=2.54E-06 Height=0.00127
MT3 3 5 4 6 Gap=0.00508 Len=0.02561 Er=9.8 Thick=2.54E-06 Height=0.00127
MT4 5 6 Wid=0.00127 Len=0.02561 Er=9.8 Thick=2.54E-06 Height=0.00127
MT5 3 5 Wid=0.00127 Len=0.00508 Er=9.8 Thick=2.54E-06 Height=0.00127
MT6 5 7 6 8 Gap=0.0002694 Len=0.02561 Er=9.8 Thick=2.54E-06 Height=0.00127
MT7 7 8 Wid=0.00127 Len=0.02561 Er=9.8 Thick=2.54E-06 Height=0.00127
MT8 7 9 8 10 Gap=0.00508 Len=0.02561 Er=9.8 Thick=2.54E-06 Height=0.00127
MT9 9 10 Wid=0.00127 Len=0.02561 Er=9.8 Thick=2.54E-06 Height=0.00127
MT10 8 10 Wid=0.00127 Len=0.00508 Er=9.8 Thick=2.54E-06 Height=0.00127
MT11 9 11 10 12 Gap=0.0008834 Len=0.02561 Er=9.8 Thick=2.54E-06 Height=0.00127
MT12 11 12 Wid=0.00127 Len=0.02561 Er=9.8 Thick=2.54E-06 Height=0.00127
MT13 11 13 12 14 Gap=0.00508 Len=0.02561 Er=9.8 Thick=2.54E-06 Height=0.00127
MT14 13 14 Wid=0.00127 Len=0.02561 Er=9.8 Thick=2.54E-06 Height=0.00127
MT15 11 13 Wid=0.00127 Len=0.00508 Er=9.8 Thick=2.54E-06 Height=0.00127
MT16 13 15 14 16 Gap=0.0008834 Len=0.02561 Er=9.8 Thick=2.54E-06 Height=0.00127
MT17 15 16 Wid=0.00127 Len=0.02561 Er=9.8 Thick=2.54E-06 Height=0.00127
MT18 15 17 16 18 Gap=0.00508 Len=0.02561 Er=9.8 Thick=2.54E-06 Height=0.00127
MT19 17 18 Wid=0.00127 Len=0.02561 Er=9.8 Thick=2.54E-06 Height=0.00127
MT20 16 18 Wid=0.00127 Len=0.00508 Er=9.8 Thick=2.54E-06 Height=0.00127
MT21 17 19 18 20 Gap=0.0002694 Len=0.02561 Er=9.8 Thick=2.54E-06 Height=0.00127
MT22 19 20 Wid=0.00127 Len=0.02561 Er=9.8 Thick=2.54E-06 Height=0.00127
MT23 19 21 20 22 Gap=0.00508 Len=0.02561 Er=9.8 Thick=2.54E-06 Height=0.00127
MT24 19 21 Wid=0.00127 Len=0.00508 Er=9.8 Thick=2.54E-06 Height=0.00127
MT25 21 23 Wid=0.00127 Len=0.01137 Er=9.8 Thick=2.54E-06 Height=0.00127
MT26 23 22 Wid=0.00127 Len=0.01424 Er=9.8 Thick=2.54E-06 Height=0.00127
Rl 23 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(Rl) -160 0
.PLOT AC VP(Rl) -200 200
.PLOT AC VG(Rl) -3E-08 3E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(Rl) -0.05 0.04
.END
