*
*Length Units: Meters
*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
Rg 1 2 50
MXTcoup0 2 5 6 3 Wid=0.0009605 Gap=0.00045 Len=0.02903 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT0 4 5 Wid=0.0009605 Len=0.02903 Er=9.8 Thick=2.54E-06 Height=0.00127 Rho=1.43 Tand=0.0005
MXTcoup1 6 9 10 7 Wid=0.0006633 Gap=0.0001582 Len=0.02955 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT1 8 9 Wid=0.0006633 Len=0.02955 Er=9.8 Thick=2.54E-06 Height=0.00127 Rho=1.43 Tand=0.0005
MXTcoup2 10 13 14 11 Wid=0.0005798 Gap=0.0001159 Len=0.02969 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT2 12 13 Wid=0.0005798 Len=0.02969 Er=9.8 Thick=2.54E-06 Height=0.00127 Rho=1.43 Tand=0.0005
MXTcoup3 14 17 18 15 Wid=0.0006633 Gap=0.0001582 Len=0.02955 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT3 16 17 Wid=0.0006633 Len=0.02955 Er=9.8 Thick=2.54E-06 Height=0.00127 Rho=1.43 Tand=0.0005
MXTcoup4 18 21 22 19 Wid=0.0009605 Gap=0.00045 Len=0.02903 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT4 20 21 Wid=0.0009605 Len=0.02903 Er=9.8 Thick=2.54E-06 Height=0.00127 Rho=1.43 Tand=0.0005
Rl 22 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(Rl) -120 0
.PLOT AC VP(Rl) -200 200
.PLOT AC VG(Rl) -2E-07 5E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(Rl) -0.1 0.6
.END
