*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
L2 2 3 8.17E-09
L3 3 4 8.595E-09
C3 4 0 2.366E-12
L4 3 5 8.123E-09
L5 5 6 4.129E-09
C5 6 0 2.523E-12
L6 5 7 1.459E-09
R7 7 0 50
C9 2 8 7.438E-13
L10 8 0 1.071E-08
C11 8 9 1.496E-12
C8 2 9 1.574E-12
C13 9 10 1.287E-12
L14 10 0 1.004E-08
C15 10 11 3.582E-12
C12 9 11 3.642E-12
R16 11 0 50
*
* Compensation Elements
*
L1 2 12 2.28E-07
C1 12 0 1.111E-13
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(7) VDB(11) -200 0
.PLOT AC VP(7) VP(11) -200 200
.PLOT AC VG(7) VG(11) 0 1.8E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(7) V(11) -0.2 0.7
.END
