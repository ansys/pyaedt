*
*Length Units: Meters
*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
Rg 1 2 50
MT1 2 3 Wid=0.00127 Len=0.007534 Er=9.8 Thick=2.54E-06 Height=0.00127
MT2 2 4 Wid=0.00127 Len=0.006381 Er=9.8 Thick=2.54E-06 Height=0.00127
MT3 4 5 Wid=0.00127 Len=0.002 Er=9.8 Thick=2.54E-06 Height=0.00127
MT4 3 6 4 7 Gap=0.01391 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT5 6 7 Wid=0.00127 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT6 3 6 Wid=0.00127 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT7 6 8 7 9 Gap=7.937E-05 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT8 8 9 Wid=0.00127 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT9 8 10 9 11 Gap=0.01391 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT10 10 11 Wid=0.00127 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT11 9 11 Wid=0.00127 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT12 10 12 11 13 Gap=0.0005276 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT13 12 13 Wid=0.00127 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT14 12 14 13 15 Gap=0.01391 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT15 14 15 Wid=0.00127 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT16 12 14 Wid=0.00127 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT17 14 16 15 17 Gap=0.0005276 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT18 16 17 Wid=0.00127 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT19 16 18 17 19 Gap=0.01391 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT20 18 19 Wid=0.00127 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT21 17 19 Wid=0.00127 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT22 18 20 19 21 Gap=7.937E-05 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT23 20 21 Wid=0.00127 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT24 20 22 21 23 Gap=0.01391 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT25 20 22 Wid=0.00127 Len=0.01391 Er=9.8 Thick=2.54E-06 Height=0.00127
MT26 22 24 Wid=0.00127 Len=0.007534 Er=9.8 Thick=2.54E-06 Height=0.00127
MT27 24 23 Wid=0.00127 Len=0.006381 Er=9.8 Thick=2.54E-06 Height=0.00127
MT28 23 25 Wid=0.00127 Len=0.002 Er=9.8 Thick=2.54E-06 Height=0.00127
Rl 24 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(Rl) -140 0
.PLOT AC VP(Rl) -200 200
.PLOT AC VG(Rl) -5E-09 1.5E-08
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(Rl) -0.05 0.04
.END
