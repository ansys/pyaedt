*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
*
* Dummy Resistors Required For Spice
* Have Been Added to Net List.
*
C2 2 3 7.12E-12
C3 3 0 3.873E-12
C4 3 4 1.233E-11
Rq4 3 4 5E+10
L1 2 4 4.424E-09
C6 4 5 3.916E-12
Rq6 4 5 5E+10
C7 5 0 9.429E-12
C8 5 6 4.684E-12
Rq8 5 6 5E+10
L5 4 6 8.388E-09
R9 6 0 50
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(6) -70 0
.PLOT AC VP(6) -200 200
.PLOT AC VG(6) 0 2.5E-09
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(6) 0 0.6
.END
