*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 50
L2 2 3 3.998E-08
C2 3 0 1.737E-11
C3 2 4 4.12E-12
L4 4 5 2.459E-08
L5 5 0 9.393E-09
C6 5 0 1.079E-11
C7 5 6 4.607E-12
L8 6 7 2.199E-08
L9 7 0 1.779E-08
C10 7 0 5.694E-12
C11 7 8 2.06E-11
L12 8 9 4.918E-09
R13 9 0 50
L14 2 10 1.458E-09
C14 10 0 6.335E-13
C15 2 11 1.03E-12
L16 11 12 6.148E-09
L17 12 0 2.348E-09
C18 12 0 2.697E-12
C19 12 13 1.152E-12
L20 13 14 5.499E-09
L21 14 0 4.449E-09
C22 14 0 1.424E-12
C23 14 15 5.15E-12
L24 15 16 1.23E-09
R25 16 0 50
*
* Compensation Elements
*
L1 2 17 2.885E-08
C1 17 0 8.78E-13
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(9) VDB(16) -200 0
.PLOT AC VP(9) VP(16) -200 200
.PLOT AC VG(9) VG(16) -1E-09 8E-09
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(9) V(16) -0.2 0.7
.END
