*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
R0 1 2 {TABLE(F, 1E+08, 1, 1E+09, 1, 1E+10, 1) + J*TABLE(F, 1E+08, 0, 1E+09, 0, 1E+10, 0)}
C1 2 0 9.836E-11
L2 2 3 2.575E-10
C3 3 0 3.183E-10
L4 3 4 2.575E-10
C5 4 0 9.836E-11
R6 4 0 {TABLE(F, 1E+08, 1, 1E+09, 1, 1E+10, 1) + J*TABLE(F, 1E+08, 0, 1E+09, 0, 1E+10, 0)}
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(4) -80 0
.PLOT AC VP(4) -200 200
.PLOT AC VG(4) 0 9E-10
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(4) 0 0.6
.END
