*
*Length Units: Meters
*
V1 1 0 AC 1 PULSE 0 1 0 1.592E-13 0
Rg 1 2 50
MTSeg0 2 3 Wid=0.0007792 Len=0.01449 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT1S1 3 0 Wid=0.0007792 Len=0.018 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MTSeg1 3 4 Wid=0.0007792 Len=0.01449 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MXTcoup2 0 4 5 0 Wid=0.0003763 Gap=0.0005407 Len=0.02947 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MXTcoup3 0 5 6 0 Wid=0.0004225 Gap=0.001121 Len=0.02926 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MXTcoup4 0 6 7 0 Wid=0.0004225 Gap=0.001121 Len=0.02926 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MXTcoup5 0 7 8 0 Wid=0.0003763 Gap=0.0005407 Len=0.02947 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MTSeg6 8 9 Wid=0.0007792 Len=0.01449 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MT1S7 9 0 Wid=0.0007792 Len=0.018 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
MTSeg7 9 10 Wid=0.0007792 Len=0.01449 Er=9.8 Height=0.00127 Thick=2.54E-06 Rho=1.43 Tand=0.0005
Rl 10 0 50
*
* The Following Dummy Resistors May Be Required For Spice.
*
Rseg8 3 0 5E+09
Rseg9 4 0 5E+09
Rseg10 9 0 5E+09
*
* End Dummy Resistors
*
*
.AC DEC 200 2E+08 5E+09
.PLOT AC VDB(Rl) -180 0
.PLOT AC VP(Rl) -200 200
.PLOT AC VG(Rl) -5E-08 1.5E-07
.TRAN  5E-11 1E-08 0
.PLOT TRAN V(Rl) -0.04 0.04
.END
